// `define VIVADO

// `define M0_LED
// `define M0_SEG7
// `define M0_TIMER
`define M0_UART
